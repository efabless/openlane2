module spm (clk,
    p,
    rst,
    y,
    x);
 input clk;
 output p;
 input rst;
 input y;
 input [31:0] x;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire \csa0.hsum2 ;
 wire \csa0.sc ;
 wire \csa0.y ;
 wire \genblk1[10].csa.hsum2 ;
 wire \genblk1[10].csa.sc ;
 wire \genblk1[10].csa.sum ;
 wire \genblk1[10].csa.y ;
 wire \genblk1[11].csa.hsum2 ;
 wire \genblk1[11].csa.sc ;
 wire \genblk1[11].csa.y ;
 wire \genblk1[12].csa.hsum2 ;
 wire \genblk1[12].csa.sc ;
 wire \genblk1[12].csa.y ;
 wire \genblk1[13].csa.hsum2 ;
 wire \genblk1[13].csa.sc ;
 wire \genblk1[13].csa.y ;
 wire \genblk1[14].csa.hsum2 ;
 wire \genblk1[14].csa.sc ;
 wire \genblk1[14].csa.y ;
 wire \genblk1[15].csa.hsum2 ;
 wire \genblk1[15].csa.sc ;
 wire \genblk1[15].csa.y ;
 wire \genblk1[16].csa.hsum2 ;
 wire \genblk1[16].csa.sc ;
 wire \genblk1[16].csa.y ;
 wire \genblk1[17].csa.hsum2 ;
 wire \genblk1[17].csa.sc ;
 wire \genblk1[17].csa.y ;
 wire \genblk1[18].csa.hsum2 ;
 wire \genblk1[18].csa.sc ;
 wire \genblk1[18].csa.y ;
 wire \genblk1[19].csa.hsum2 ;
 wire \genblk1[19].csa.sc ;
 wire \genblk1[19].csa.y ;
 wire \genblk1[1].csa.hsum2 ;
 wire \genblk1[1].csa.sc ;
 wire \genblk1[1].csa.y ;
 wire \genblk1[20].csa.hsum2 ;
 wire \genblk1[20].csa.sc ;
 wire \genblk1[20].csa.y ;
 wire \genblk1[21].csa.hsum2 ;
 wire \genblk1[21].csa.sc ;
 wire \genblk1[21].csa.y ;
 wire \genblk1[22].csa.hsum2 ;
 wire \genblk1[22].csa.sc ;
 wire \genblk1[22].csa.y ;
 wire \genblk1[23].csa.hsum2 ;
 wire \genblk1[23].csa.sc ;
 wire \genblk1[23].csa.y ;
 wire \genblk1[24].csa.hsum2 ;
 wire \genblk1[24].csa.sc ;
 wire \genblk1[24].csa.y ;
 wire \genblk1[25].csa.hsum2 ;
 wire \genblk1[25].csa.sc ;
 wire \genblk1[25].csa.y ;
 wire \genblk1[26].csa.hsum2 ;
 wire \genblk1[26].csa.sc ;
 wire \genblk1[26].csa.y ;
 wire \genblk1[27].csa.hsum2 ;
 wire \genblk1[27].csa.sc ;
 wire \genblk1[27].csa.y ;
 wire \genblk1[28].csa.hsum2 ;
 wire \genblk1[28].csa.sc ;
 wire \genblk1[28].csa.y ;
 wire \genblk1[29].csa.hsum2 ;
 wire \genblk1[29].csa.sc ;
 wire \genblk1[29].csa.y ;
 wire \genblk1[2].csa.hsum2 ;
 wire \genblk1[2].csa.sc ;
 wire \genblk1[2].csa.y ;
 wire \genblk1[30].csa.hsum2 ;
 wire \genblk1[30].csa.sc ;
 wire \genblk1[30].csa.y ;
 wire \genblk1[3].csa.hsum2 ;
 wire \genblk1[3].csa.sc ;
 wire \genblk1[3].csa.y ;
 wire \genblk1[4].csa.hsum2 ;
 wire \genblk1[4].csa.sc ;
 wire \genblk1[4].csa.y ;
 wire \genblk1[5].csa.hsum2 ;
 wire \genblk1[5].csa.sc ;
 wire \genblk1[5].csa.y ;
 wire \genblk1[6].csa.hsum2 ;
 wire \genblk1[6].csa.sc ;
 wire \genblk1[6].csa.y ;
 wire \genblk1[7].csa.hsum2 ;
 wire \genblk1[7].csa.sc ;
 wire \genblk1[7].csa.y ;
 wire \genblk1[8].csa.hsum2 ;
 wire \genblk1[8].csa.sc ;
 wire \genblk1[8].csa.y ;
 wire \genblk1[9].csa.hsum2 ;
 wire \genblk1[9].csa.sc ;
 wire \tcmp.z ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;

 sky130_fd_sc_hd__xor2_1 _192_ (.A(\csa0.sc ),
    .B(\csa0.y ),
    .X(_097_));
 sky130_fd_sc_hd__and2_1 _193_ (.A(\csa0.sc ),
    .B(\csa0.y ),
    .X(_098_));
 sky130_fd_sc_hd__a31o_1 _194_ (.A1(net36),
    .A2(net2),
    .A3(_097_),
    .B1(_098_),
    .X(_000_));
 sky130_fd_sc_hd__nand2_1 _195_ (.A(net36),
    .B(net2),
    .Y(_099_));
 sky130_fd_sc_hd__xnor2_1 _196_ (.A(_099_),
    .B(_097_),
    .Y(\csa0.hsum2 ));
 sky130_fd_sc_hd__a21o_1 _197_ (.A1(net41),
    .A2(net26),
    .B1(\tcmp.z ),
    .X(_032_));
 sky130_fd_sc_hd__nand3_1 _198_ (.A(net41),
    .B(net26),
    .C(\tcmp.z ),
    .Y(_100_));
 sky130_fd_sc_hd__and2_1 _199_ (.A(_032_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(_101_),
    .X(_031_));
 sky130_fd_sc_hd__xor2_1 _201_ (.A(\genblk1[1].csa.sc ),
    .B(\genblk1[1].csa.y ),
    .X(_102_));
 sky130_fd_sc_hd__and2_1 _202_ (.A(\genblk1[1].csa.sc ),
    .B(\genblk1[1].csa.y ),
    .X(_103_));
 sky130_fd_sc_hd__a31o_1 _203_ (.A1(net36),
    .A2(net13),
    .A3(_102_),
    .B1(_103_),
    .X(_011_));
 sky130_fd_sc_hd__nand2_1 _204_ (.A(net36),
    .B(net13),
    .Y(_104_));
 sky130_fd_sc_hd__xnor2_1 _205_ (.A(_104_),
    .B(_102_),
    .Y(\genblk1[1].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _206_ (.A(\genblk1[2].csa.sc ),
    .B(\genblk1[2].csa.y ),
    .X(_105_));
 sky130_fd_sc_hd__and2_1 _207_ (.A(\genblk1[2].csa.sc ),
    .B(\genblk1[2].csa.y ),
    .X(_106_));
 sky130_fd_sc_hd__a31o_1 _208_ (.A1(net37),
    .A2(net24),
    .A3(_105_),
    .B1(_106_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_1 _209_ (.A(net36),
    .B(net24),
    .Y(_107_));
 sky130_fd_sc_hd__xnor2_1 _210_ (.A(_107_),
    .B(_105_),
    .Y(\genblk1[2].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _211_ (.A(\genblk1[3].csa.sc ),
    .B(\genblk1[3].csa.y ),
    .X(_108_));
 sky130_fd_sc_hd__and2_1 _212_ (.A(\genblk1[3].csa.sc ),
    .B(\genblk1[3].csa.y ),
    .X(_109_));
 sky130_fd_sc_hd__a31o_1 _213_ (.A1(net37),
    .A2(net27),
    .A3(_108_),
    .B1(_109_),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _214_ (.A(net37),
    .B(net27),
    .Y(_110_));
 sky130_fd_sc_hd__xnor2_1 _215_ (.A(_110_),
    .B(_108_),
    .Y(\genblk1[3].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _216_ (.A(\genblk1[4].csa.sc ),
    .B(\genblk1[4].csa.y ),
    .X(_111_));
 sky130_fd_sc_hd__and2_1 _217_ (.A(\genblk1[4].csa.sc ),
    .B(\genblk1[4].csa.y ),
    .X(_112_));
 sky130_fd_sc_hd__a31o_1 _218_ (.A1(net37),
    .A2(net28),
    .A3(_111_),
    .B1(_112_),
    .X(_025_));
 sky130_fd_sc_hd__nand2_1 _219_ (.A(net37),
    .B(net28),
    .Y(_113_));
 sky130_fd_sc_hd__xnor2_1 _220_ (.A(_113_),
    .B(_111_),
    .Y(\genblk1[4].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _221_ (.A(\genblk1[5].csa.sc ),
    .B(\genblk1[5].csa.y ),
    .X(_114_));
 sky130_fd_sc_hd__and2_1 _222_ (.A(\genblk1[5].csa.sc ),
    .B(\genblk1[5].csa.y ),
    .X(_115_));
 sky130_fd_sc_hd__a31o_1 _223_ (.A1(net37),
    .A2(net29),
    .A3(_114_),
    .B1(_115_),
    .X(_026_));
 sky130_fd_sc_hd__nand2_1 _224_ (.A(net37),
    .B(net29),
    .Y(_116_));
 sky130_fd_sc_hd__xnor2_1 _225_ (.A(_116_),
    .B(_114_),
    .Y(\genblk1[5].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _226_ (.A(\genblk1[6].csa.sc ),
    .B(\genblk1[6].csa.y ),
    .X(_117_));
 sky130_fd_sc_hd__and2_1 _227_ (.A(\genblk1[6].csa.sc ),
    .B(\genblk1[6].csa.y ),
    .X(_118_));
 sky130_fd_sc_hd__a31o_1 _228_ (.A1(net37),
    .A2(net30),
    .A3(_117_),
    .B1(_118_),
    .X(_027_));
 sky130_fd_sc_hd__nand2_1 _229_ (.A(net37),
    .B(net30),
    .Y(_119_));
 sky130_fd_sc_hd__xnor2_1 _230_ (.A(_119_),
    .B(_117_),
    .Y(\genblk1[6].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _231_ (.A(\genblk1[7].csa.sc ),
    .B(\genblk1[7].csa.y ),
    .X(_120_));
 sky130_fd_sc_hd__and2_1 _232_ (.A(\genblk1[7].csa.sc ),
    .B(\genblk1[7].csa.y ),
    .X(_121_));
 sky130_fd_sc_hd__a31o_1 _233_ (.A1(net36),
    .A2(net31),
    .A3(_120_),
    .B1(_121_),
    .X(_028_));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(net36),
    .B(net31),
    .Y(_122_));
 sky130_fd_sc_hd__xnor2_1 _235_ (.A(_122_),
    .B(_120_),
    .Y(\genblk1[7].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _236_ (.A(\genblk1[8].csa.sc ),
    .B(\genblk1[8].csa.y ),
    .X(_123_));
 sky130_fd_sc_hd__and2_1 _237_ (.A(\genblk1[8].csa.sc ),
    .B(\genblk1[8].csa.y ),
    .X(_124_));
 sky130_fd_sc_hd__a31o_1 _238_ (.A1(net36),
    .A2(net32),
    .A3(_123_),
    .B1(_124_),
    .X(_029_));
 sky130_fd_sc_hd__nand2_1 _239_ (.A(net36),
    .B(net32),
    .Y(_125_));
 sky130_fd_sc_hd__xnor2_1 _240_ (.A(_125_),
    .B(_123_),
    .Y(\genblk1[8].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _241_ (.A(\genblk1[9].csa.sc ),
    .B(\genblk1[10].csa.sum ),
    .X(_126_));
 sky130_fd_sc_hd__and2_1 _242_ (.A(\genblk1[9].csa.sc ),
    .B(\genblk1[10].csa.sum ),
    .X(_127_));
 sky130_fd_sc_hd__a31o_1 _243_ (.A1(net36),
    .A2(net33),
    .A3(_126_),
    .B1(_127_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _244_ (.A(net38),
    .B(net33),
    .Y(_128_));
 sky130_fd_sc_hd__xnor2_1 _245_ (.A(_128_),
    .B(_126_),
    .Y(\genblk1[9].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _246_ (.A(\genblk1[10].csa.sc ),
    .B(\genblk1[10].csa.y ),
    .X(_129_));
 sky130_fd_sc_hd__and2_1 _247_ (.A(\genblk1[10].csa.sc ),
    .B(\genblk1[10].csa.y ),
    .X(_130_));
 sky130_fd_sc_hd__a31o_1 _248_ (.A1(net38),
    .A2(net3),
    .A3(_129_),
    .B1(_130_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(net38),
    .B(net3),
    .Y(_131_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_131_),
    .B(_129_),
    .Y(\genblk1[10].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _251_ (.A(\genblk1[11].csa.sc ),
    .B(\genblk1[11].csa.y ),
    .X(_132_));
 sky130_fd_sc_hd__and2_1 _252_ (.A(\genblk1[11].csa.sc ),
    .B(\genblk1[11].csa.y ),
    .X(_133_));
 sky130_fd_sc_hd__a31o_1 _253_ (.A1(net37),
    .A2(net4),
    .A3(_132_),
    .B1(_133_),
    .X(_002_));
 sky130_fd_sc_hd__nand2_1 _254_ (.A(net38),
    .B(net4),
    .Y(_134_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_134_),
    .B(_132_),
    .Y(\genblk1[11].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _256_ (.A(\genblk1[12].csa.sc ),
    .B(\genblk1[12].csa.y ),
    .X(_135_));
 sky130_fd_sc_hd__and2_1 _257_ (.A(\genblk1[12].csa.sc ),
    .B(\genblk1[12].csa.y ),
    .X(_136_));
 sky130_fd_sc_hd__a31o_1 _258_ (.A1(net38),
    .A2(net5),
    .A3(_135_),
    .B1(_136_),
    .X(_003_));
 sky130_fd_sc_hd__nand2_1 _259_ (.A(net38),
    .B(net5),
    .Y(_137_));
 sky130_fd_sc_hd__xnor2_1 _260_ (.A(_137_),
    .B(_135_),
    .Y(\genblk1[12].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _261_ (.A(\genblk1[13].csa.sc ),
    .B(\genblk1[13].csa.y ),
    .X(_138_));
 sky130_fd_sc_hd__and2_1 _262_ (.A(\genblk1[13].csa.sc ),
    .B(\genblk1[13].csa.y ),
    .X(_139_));
 sky130_fd_sc_hd__a31o_1 _263_ (.A1(net38),
    .A2(net6),
    .A3(_138_),
    .B1(_139_),
    .X(_004_));
 sky130_fd_sc_hd__nand2_1 _264_ (.A(net38),
    .B(net6),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_1 _265_ (.A(_140_),
    .B(_138_),
    .Y(\genblk1[13].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _266_ (.A(\genblk1[14].csa.sc ),
    .B(\genblk1[14].csa.y ),
    .X(_141_));
 sky130_fd_sc_hd__and2_1 _267_ (.A(\genblk1[14].csa.sc ),
    .B(\genblk1[14].csa.y ),
    .X(_142_));
 sky130_fd_sc_hd__a31o_1 _268_ (.A1(net41),
    .A2(net7),
    .A3(_141_),
    .B1(_142_),
    .X(_005_));
 sky130_fd_sc_hd__nand2_1 _269_ (.A(net41),
    .B(net7),
    .Y(_143_));
 sky130_fd_sc_hd__xnor2_1 _270_ (.A(_143_),
    .B(_141_),
    .Y(\genblk1[14].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _271_ (.A(\genblk1[15].csa.sc ),
    .B(\genblk1[15].csa.y ),
    .X(_144_));
 sky130_fd_sc_hd__and2_1 _272_ (.A(\genblk1[15].csa.sc ),
    .B(\genblk1[15].csa.y ),
    .X(_145_));
 sky130_fd_sc_hd__a31o_1 _273_ (.A1(net41),
    .A2(net8),
    .A3(_144_),
    .B1(_145_),
    .X(_006_));
 sky130_fd_sc_hd__nand2_1 _274_ (.A(net41),
    .B(net8),
    .Y(_146_));
 sky130_fd_sc_hd__xnor2_1 _275_ (.A(_146_),
    .B(_144_),
    .Y(\genblk1[15].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _276_ (.A(\genblk1[16].csa.sc ),
    .B(\genblk1[16].csa.y ),
    .X(_147_));
 sky130_fd_sc_hd__and2_1 _277_ (.A(\genblk1[16].csa.sc ),
    .B(\genblk1[16].csa.y ),
    .X(_148_));
 sky130_fd_sc_hd__a31o_1 _278_ (.A1(net39),
    .A2(net9),
    .A3(_147_),
    .B1(_148_),
    .X(_007_));
 sky130_fd_sc_hd__nand2_1 _279_ (.A(net39),
    .B(net9),
    .Y(_149_));
 sky130_fd_sc_hd__xnor2_1 _280_ (.A(_149_),
    .B(_147_),
    .Y(\genblk1[16].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _281_ (.A(\genblk1[17].csa.sc ),
    .B(\genblk1[17].csa.y ),
    .X(_150_));
 sky130_fd_sc_hd__and2_1 _282_ (.A(\genblk1[17].csa.sc ),
    .B(\genblk1[17].csa.y ),
    .X(_151_));
 sky130_fd_sc_hd__a31o_1 _283_ (.A1(net39),
    .A2(net10),
    .A3(_150_),
    .B1(_151_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _284_ (.A(net39),
    .B(net10),
    .Y(_152_));
 sky130_fd_sc_hd__xnor2_1 _285_ (.A(_152_),
    .B(_150_),
    .Y(\genblk1[17].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _286_ (.A(\genblk1[18].csa.sc ),
    .B(\genblk1[18].csa.y ),
    .X(_153_));
 sky130_fd_sc_hd__and2_1 _287_ (.A(\genblk1[18].csa.sc ),
    .B(\genblk1[18].csa.y ),
    .X(_154_));
 sky130_fd_sc_hd__a31o_1 _288_ (.A1(net39),
    .A2(net11),
    .A3(_153_),
    .B1(_154_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(net39),
    .B(net11),
    .Y(_155_));
 sky130_fd_sc_hd__xnor2_1 _290_ (.A(_155_),
    .B(_153_),
    .Y(\genblk1[18].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _291_ (.A(\genblk1[19].csa.sc ),
    .B(\genblk1[19].csa.y ),
    .X(_156_));
 sky130_fd_sc_hd__and2_1 _292_ (.A(\genblk1[19].csa.sc ),
    .B(\genblk1[19].csa.y ),
    .X(_157_));
 sky130_fd_sc_hd__a31o_1 _293_ (.A1(net39),
    .A2(net12),
    .A3(_156_),
    .B1(_157_),
    .X(_010_));
 sky130_fd_sc_hd__nand2_1 _294_ (.A(net39),
    .B(net12),
    .Y(_158_));
 sky130_fd_sc_hd__xnor2_1 _295_ (.A(_158_),
    .B(_156_),
    .Y(\genblk1[19].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _296_ (.A(\genblk1[20].csa.sc ),
    .B(\genblk1[20].csa.y ),
    .X(_159_));
 sky130_fd_sc_hd__and2_1 _297_ (.A(\genblk1[20].csa.sc ),
    .B(\genblk1[20].csa.y ),
    .X(_160_));
 sky130_fd_sc_hd__a31o_1 _298_ (.A1(net41),
    .A2(net14),
    .A3(_159_),
    .B1(_160_),
    .X(_012_));
 sky130_fd_sc_hd__nand2_1 _299_ (.A(net41),
    .B(net14),
    .Y(_161_));
 sky130_fd_sc_hd__xnor2_1 _300_ (.A(_161_),
    .B(_159_),
    .Y(\genblk1[20].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _301_ (.A(\genblk1[21].csa.sc ),
    .B(\genblk1[21].csa.y ),
    .X(_162_));
 sky130_fd_sc_hd__and2_1 _302_ (.A(\genblk1[21].csa.sc ),
    .B(\genblk1[21].csa.y ),
    .X(_163_));
 sky130_fd_sc_hd__a31o_1 _303_ (.A1(net41),
    .A2(net15),
    .A3(_162_),
    .B1(_163_),
    .X(_013_));
 sky130_fd_sc_hd__nand2_1 _304_ (.A(net41),
    .B(net15),
    .Y(_164_));
 sky130_fd_sc_hd__xnor2_1 _305_ (.A(_164_),
    .B(_162_),
    .Y(\genblk1[21].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _306_ (.A(\genblk1[22].csa.sc ),
    .B(\genblk1[22].csa.y ),
    .X(_165_));
 sky130_fd_sc_hd__and2_1 _307_ (.A(\genblk1[22].csa.sc ),
    .B(\genblk1[22].csa.y ),
    .X(_166_));
 sky130_fd_sc_hd__a31o_1 _308_ (.A1(net42),
    .A2(net16),
    .A3(_165_),
    .B1(_166_),
    .X(_014_));
 sky130_fd_sc_hd__nand2_1 _309_ (.A(net42),
    .B(net16),
    .Y(_167_));
 sky130_fd_sc_hd__xnor2_1 _310_ (.A(_167_),
    .B(_165_),
    .Y(\genblk1[22].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _311_ (.A(\genblk1[23].csa.sc ),
    .B(\genblk1[23].csa.y ),
    .X(_168_));
 sky130_fd_sc_hd__and2_1 _312_ (.A(\genblk1[23].csa.sc ),
    .B(\genblk1[23].csa.y ),
    .X(_169_));
 sky130_fd_sc_hd__a31o_1 _313_ (.A1(net42),
    .A2(net17),
    .A3(_168_),
    .B1(_169_),
    .X(_015_));
 sky130_fd_sc_hd__nand2_1 _314_ (.A(net42),
    .B(net17),
    .Y(_170_));
 sky130_fd_sc_hd__xnor2_1 _315_ (.A(_170_),
    .B(_168_),
    .Y(\genblk1[23].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _316_ (.A(\genblk1[24].csa.sc ),
    .B(\genblk1[24].csa.y ),
    .X(_171_));
 sky130_fd_sc_hd__and2_1 _317_ (.A(\genblk1[24].csa.sc ),
    .B(\genblk1[24].csa.y ),
    .X(_172_));
 sky130_fd_sc_hd__a31o_1 _318_ (.A1(net39),
    .A2(net18),
    .A3(_171_),
    .B1(_172_),
    .X(_016_));
 sky130_fd_sc_hd__nand2_1 _319_ (.A(net39),
    .B(net18),
    .Y(_173_));
 sky130_fd_sc_hd__xnor2_1 _320_ (.A(_173_),
    .B(_171_),
    .Y(\genblk1[24].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _321_ (.A(\genblk1[25].csa.sc ),
    .B(\genblk1[25].csa.y ),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _322_ (.A(\genblk1[25].csa.sc ),
    .B(\genblk1[25].csa.y ),
    .X(_175_));
 sky130_fd_sc_hd__a31o_1 _323_ (.A1(net40),
    .A2(net19),
    .A3(_174_),
    .B1(_175_),
    .X(_017_));
 sky130_fd_sc_hd__nand2_1 _324_ (.A(net40),
    .B(net19),
    .Y(_176_));
 sky130_fd_sc_hd__xnor2_1 _325_ (.A(_176_),
    .B(_174_),
    .Y(\genblk1[25].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _326_ (.A(\genblk1[26].csa.sc ),
    .B(\genblk1[26].csa.y ),
    .X(_177_));
 sky130_fd_sc_hd__and2_1 _327_ (.A(\genblk1[26].csa.sc ),
    .B(\genblk1[26].csa.y ),
    .X(_178_));
 sky130_fd_sc_hd__a31o_1 _328_ (.A1(net40),
    .A2(net20),
    .A3(_177_),
    .B1(_178_),
    .X(_018_));
 sky130_fd_sc_hd__nand2_1 _329_ (.A(net40),
    .B(net20),
    .Y(_179_));
 sky130_fd_sc_hd__xnor2_1 _330_ (.A(_179_),
    .B(_177_),
    .Y(\genblk1[26].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _331_ (.A(\genblk1[27].csa.sc ),
    .B(\genblk1[27].csa.y ),
    .X(_180_));
 sky130_fd_sc_hd__and2_1 _332_ (.A(\genblk1[27].csa.sc ),
    .B(\genblk1[27].csa.y ),
    .X(_181_));
 sky130_fd_sc_hd__a31o_1 _333_ (.A1(net40),
    .A2(net21),
    .A3(_180_),
    .B1(_181_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _334_ (.A(net40),
    .B(net21),
    .Y(_182_));
 sky130_fd_sc_hd__xnor2_1 _335_ (.A(_182_),
    .B(_180_),
    .Y(\genblk1[27].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _336_ (.A(\genblk1[28].csa.sc ),
    .B(\genblk1[28].csa.y ),
    .X(_183_));
 sky130_fd_sc_hd__and2_1 _337_ (.A(\genblk1[28].csa.sc ),
    .B(\genblk1[28].csa.y ),
    .X(_184_));
 sky130_fd_sc_hd__a31o_1 _338_ (.A1(net40),
    .A2(net22),
    .A3(_183_),
    .B1(_184_),
    .X(_020_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(net40),
    .B(net22),
    .Y(_185_));
 sky130_fd_sc_hd__xnor2_1 _340_ (.A(_185_),
    .B(_183_),
    .Y(\genblk1[28].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _341_ (.A(\genblk1[29].csa.sc ),
    .B(\genblk1[29].csa.y ),
    .X(_186_));
 sky130_fd_sc_hd__and2_1 _342_ (.A(\genblk1[29].csa.sc ),
    .B(\genblk1[29].csa.y ),
    .X(_187_));
 sky130_fd_sc_hd__a31o_1 _343_ (.A1(net42),
    .A2(net23),
    .A3(_186_),
    .B1(_187_),
    .X(_021_));
 sky130_fd_sc_hd__nand2_1 _344_ (.A(net42),
    .B(net23),
    .Y(_188_));
 sky130_fd_sc_hd__xnor2_1 _345_ (.A(_188_),
    .B(_186_),
    .Y(\genblk1[29].csa.hsum2 ));
 sky130_fd_sc_hd__xor2_1 _346_ (.A(\genblk1[30].csa.sc ),
    .B(\genblk1[30].csa.y ),
    .X(_189_));
 sky130_fd_sc_hd__and2_1 _347_ (.A(\genblk1[30].csa.sc ),
    .B(\genblk1[30].csa.y ),
    .X(_190_));
 sky130_fd_sc_hd__a31o_1 _348_ (.A1(net42),
    .A2(net25),
    .A3(_189_),
    .B1(_190_),
    .X(_023_));
 sky130_fd_sc_hd__nand2_1 _349_ (.A(net42),
    .B(net25),
    .Y(_191_));
 sky130_fd_sc_hd__xnor2_1 _350_ (.A(_191_),
    .B(_189_),
    .Y(\genblk1[30].csa.hsum2 ));
 sky130_fd_sc_hd__inv_2 _351_ (.A(net44),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _352_ (.A(net44),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(net49),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _354_ (.A(net49),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _355_ (.A(net44),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _356_ (.A(net44),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _357_ (.A(net46),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _358_ (.A(net44),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _359_ (.A(net46),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _360_ (.A(net46),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(net46),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _362_ (.A(net46),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _363_ (.A(net46),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _364_ (.A(net46),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _365_ (.A(net46),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _366_ (.A(net46),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _367_ (.A(net44),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _368_ (.A(net46),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _369_ (.A(net44),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _370_ (.A(net44),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net44),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _372_ (.A(net44),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _373_ (.A(net45),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _374_ (.A(net45),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(net47),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _376_ (.A(net45),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(net47),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _378_ (.A(net47),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _379_ (.A(net47),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(net47),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(net47),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(net50),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(net47),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(net50),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _385_ (.A(net45),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _386_ (.A(net48),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(net45),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net45),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net48),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net48),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(net48),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(net48),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(net50),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(net50),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(net50),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(net50),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(net49),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(net49),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(net49),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(net49),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(net48),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(net49),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _403_ (.A(net48),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(net48),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(net48),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _406_ (.A(net48),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(net51),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(net51),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(net51),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _410_ (.A(net51),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(net49),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _412_ (.A(net49),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _413_ (.A(net50),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _414_ (.A(net49),
    .Y(_096_));
 sky130_fd_sc_hd__dfrtp_1 _415_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_033_),
    .Q(\csa0.sc ));
 sky130_fd_sc_hd__dfrtp_1 _416_ (.CLK(clk),
    .D(\csa0.hsum2 ),
    .RESET_B(_034_),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _417_ (.CLK(clk),
    .D(_032_),
    .RESET_B(_035_),
    .Q(\tcmp.z ));
 sky130_fd_sc_hd__dfrtp_1 _418_ (.CLK(clk),
    .D(_031_),
    .RESET_B(_036_),
    .Q(\genblk1[30].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _419_ (.CLK(clk),
    .D(_011_),
    .RESET_B(_037_),
    .Q(\genblk1[1].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _420_ (.CLK(clk),
    .D(\genblk1[1].csa.hsum2 ),
    .RESET_B(_038_),
    .Q(\csa0.y ));
 sky130_fd_sc_hd__dfrtp_1 _421_ (.CLK(clk),
    .D(_022_),
    .RESET_B(_039_),
    .Q(\genblk1[2].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _422_ (.CLK(clk),
    .D(\genblk1[2].csa.hsum2 ),
    .RESET_B(_040_),
    .Q(\genblk1[1].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _423_ (.CLK(clk),
    .D(_024_),
    .RESET_B(_041_),
    .Q(\genblk1[3].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _424_ (.CLK(clk),
    .D(\genblk1[3].csa.hsum2 ),
    .RESET_B(_042_),
    .Q(\genblk1[2].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _425_ (.CLK(clk),
    .D(_025_),
    .RESET_B(_043_),
    .Q(\genblk1[4].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _426_ (.CLK(clk),
    .D(\genblk1[4].csa.hsum2 ),
    .RESET_B(_044_),
    .Q(\genblk1[3].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _427_ (.CLK(clk),
    .D(_026_),
    .RESET_B(_045_),
    .Q(\genblk1[5].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _428_ (.CLK(clk),
    .D(\genblk1[5].csa.hsum2 ),
    .RESET_B(_046_),
    .Q(\genblk1[4].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _429_ (.CLK(clk),
    .D(_027_),
    .RESET_B(_047_),
    .Q(\genblk1[6].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _430_ (.CLK(clk),
    .D(\genblk1[6].csa.hsum2 ),
    .RESET_B(_048_),
    .Q(\genblk1[5].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _431_ (.CLK(clk),
    .D(_028_),
    .RESET_B(_049_),
    .Q(\genblk1[7].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _432_ (.CLK(clk),
    .D(\genblk1[7].csa.hsum2 ),
    .RESET_B(_050_),
    .Q(\genblk1[6].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _433_ (.CLK(clk),
    .D(_029_),
    .RESET_B(_051_),
    .Q(\genblk1[8].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _434_ (.CLK(clk),
    .D(\genblk1[8].csa.hsum2 ),
    .RESET_B(_052_),
    .Q(\genblk1[7].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _435_ (.CLK(clk),
    .D(_030_),
    .RESET_B(_053_),
    .Q(\genblk1[9].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _436_ (.CLK(clk),
    .D(\genblk1[9].csa.hsum2 ),
    .RESET_B(_054_),
    .Q(\genblk1[8].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _437_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_055_),
    .Q(\genblk1[10].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _438_ (.CLK(clk),
    .D(\genblk1[10].csa.hsum2 ),
    .RESET_B(_056_),
    .Q(\genblk1[10].csa.sum ));
 sky130_fd_sc_hd__dfrtp_1 _439_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_057_),
    .Q(\genblk1[11].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _440_ (.CLK(clk),
    .D(\genblk1[11].csa.hsum2 ),
    .RESET_B(_058_),
    .Q(\genblk1[10].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _441_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_059_),
    .Q(\genblk1[12].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _442_ (.CLK(clk),
    .D(\genblk1[12].csa.hsum2 ),
    .RESET_B(_060_),
    .Q(\genblk1[11].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _443_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_061_),
    .Q(\genblk1[13].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _444_ (.CLK(clk),
    .D(\genblk1[13].csa.hsum2 ),
    .RESET_B(_062_),
    .Q(\genblk1[12].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _445_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_063_),
    .Q(\genblk1[14].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _446_ (.CLK(clk),
    .D(\genblk1[14].csa.hsum2 ),
    .RESET_B(_064_),
    .Q(\genblk1[13].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _447_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_065_),
    .Q(\genblk1[15].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _448_ (.CLK(clk),
    .D(\genblk1[15].csa.hsum2 ),
    .RESET_B(_066_),
    .Q(\genblk1[14].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _449_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_067_),
    .Q(\genblk1[16].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _450_ (.CLK(clk),
    .D(\genblk1[16].csa.hsum2 ),
    .RESET_B(_068_),
    .Q(\genblk1[15].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _451_ (.CLK(clk),
    .D(_008_),
    .RESET_B(_069_),
    .Q(\genblk1[17].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _452_ (.CLK(clk),
    .D(\genblk1[17].csa.hsum2 ),
    .RESET_B(_070_),
    .Q(\genblk1[16].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _453_ (.CLK(clk),
    .D(_009_),
    .RESET_B(_071_),
    .Q(\genblk1[18].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _454_ (.CLK(clk),
    .D(\genblk1[18].csa.hsum2 ),
    .RESET_B(_072_),
    .Q(\genblk1[17].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _455_ (.CLK(clk),
    .D(_010_),
    .RESET_B(_073_),
    .Q(\genblk1[19].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _456_ (.CLK(clk),
    .D(\genblk1[19].csa.hsum2 ),
    .RESET_B(_074_),
    .Q(\genblk1[18].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _457_ (.CLK(clk),
    .D(_012_),
    .RESET_B(_075_),
    .Q(\genblk1[20].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _458_ (.CLK(clk),
    .D(\genblk1[20].csa.hsum2 ),
    .RESET_B(_076_),
    .Q(\genblk1[19].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _459_ (.CLK(clk),
    .D(_013_),
    .RESET_B(_077_),
    .Q(\genblk1[21].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _460_ (.CLK(clk),
    .D(\genblk1[21].csa.hsum2 ),
    .RESET_B(_078_),
    .Q(\genblk1[20].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _461_ (.CLK(clk),
    .D(_014_),
    .RESET_B(_079_),
    .Q(\genblk1[22].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _462_ (.CLK(clk),
    .D(\genblk1[22].csa.hsum2 ),
    .RESET_B(_080_),
    .Q(\genblk1[21].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _463_ (.CLK(clk),
    .D(_015_),
    .RESET_B(_081_),
    .Q(\genblk1[23].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(clk),
    .D(\genblk1[23].csa.hsum2 ),
    .RESET_B(_082_),
    .Q(\genblk1[22].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(clk),
    .D(_016_),
    .RESET_B(_083_),
    .Q(\genblk1[24].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(clk),
    .D(\genblk1[24].csa.hsum2 ),
    .RESET_B(_084_),
    .Q(\genblk1[23].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _467_ (.CLK(clk),
    .D(_017_),
    .RESET_B(_085_),
    .Q(\genblk1[25].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _468_ (.CLK(clk),
    .D(\genblk1[25].csa.hsum2 ),
    .RESET_B(_086_),
    .Q(\genblk1[24].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _469_ (.CLK(clk),
    .D(_018_),
    .RESET_B(_087_),
    .Q(\genblk1[26].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _470_ (.CLK(clk),
    .D(\genblk1[26].csa.hsum2 ),
    .RESET_B(_088_),
    .Q(\genblk1[25].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _471_ (.CLK(clk),
    .D(_019_),
    .RESET_B(_089_),
    .Q(\genblk1[27].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _472_ (.CLK(clk),
    .D(\genblk1[27].csa.hsum2 ),
    .RESET_B(_090_),
    .Q(\genblk1[26].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _473_ (.CLK(clk),
    .D(_020_),
    .RESET_B(_091_),
    .Q(\genblk1[28].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _474_ (.CLK(clk),
    .D(\genblk1[28].csa.hsum2 ),
    .RESET_B(_092_),
    .Q(\genblk1[27].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _475_ (.CLK(clk),
    .D(_021_),
    .RESET_B(_093_),
    .Q(\genblk1[29].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(clk),
    .D(\genblk1[29].csa.hsum2 ),
    .RESET_B(_094_),
    .Q(\genblk1[28].csa.y ));
 sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(clk),
    .D(_023_),
    .RESET_B(_095_),
    .Q(\genblk1[30].csa.sc ));
 sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(clk),
    .D(\genblk1[30].csa.hsum2 ),
    .RESET_B(_096_),
    .Q(\genblk1[29].csa.y ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(x[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(x[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(x[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(x[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(x[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(x[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(x[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(x[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(x[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(x[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(x[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(x[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(x[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(x[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(x[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(x[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(x[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(x[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(x[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(x[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(x[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(x[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(x[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(x[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(x[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(x[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(x[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(x[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(x[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(x[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(x[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(x[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(y),
    .X(net34));
 sky130_fd_sc_hd__buf_6 output35 (.A(net35),
    .X(p));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net43),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net43),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net43),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net34),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net52),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net52),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(net52),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net52),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net51),
    .X(net48));
 sky130_fd_sc_hd__buf_4 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net1),
    .X(net52));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_188 ();
endmodule
